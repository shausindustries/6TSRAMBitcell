magic
tech sky130A
timestamp 1770843875
<< nwell >>
rect -75 -35 245 200
<< nmos >>
rect -115 -180 -100 -120
rect 0 -180 15 -120
rect 165 -180 180 -120
rect 280 -180 295 -120
<< pmos >>
rect 0 -15 15 80
rect 165 -15 180 80
<< ndiff >>
rect -150 -130 -115 -120
rect -150 -170 -145 -130
rect -125 -170 -115 -130
rect -150 -180 -115 -170
rect -100 -130 -65 -120
rect -100 -170 -90 -130
rect -70 -170 -65 -130
rect -100 -180 -65 -170
rect -35 -130 0 -120
rect -35 -170 -30 -130
rect -10 -170 0 -130
rect -35 -180 0 -170
rect 15 -130 50 -120
rect 15 -170 25 -130
rect 45 -170 50 -130
rect 15 -180 50 -170
rect 130 -130 165 -120
rect 130 -170 135 -130
rect 155 -170 165 -130
rect 130 -180 165 -170
rect 180 -130 215 -120
rect 180 -170 190 -130
rect 210 -170 215 -130
rect 180 -180 215 -170
rect 245 -130 280 -120
rect 245 -170 250 -130
rect 270 -170 280 -130
rect 245 -180 280 -170
rect 295 -130 330 -120
rect 295 -170 305 -130
rect 325 -170 330 -130
rect 295 -180 330 -170
<< pdiff >>
rect -40 65 0 80
rect -40 0 -30 65
rect -10 0 0 65
rect -40 -15 0 0
rect 15 65 55 80
rect 15 0 25 65
rect 45 0 55 65
rect 15 -15 55 0
rect 125 65 165 80
rect 125 0 135 65
rect 155 0 165 65
rect 125 -15 165 0
rect 180 65 220 80
rect 180 0 190 65
rect 210 0 220 65
rect 180 -15 220 0
<< ndiffc >>
rect -145 -170 -125 -130
rect -90 -170 -70 -130
rect -30 -170 -10 -130
rect 25 -170 45 -130
rect 135 -170 155 -130
rect 190 -170 210 -130
rect 250 -170 270 -130
rect 305 -170 325 -130
<< pdiffc >>
rect -30 0 -10 65
rect 25 0 45 65
rect 135 0 155 65
rect 190 0 210 65
<< psubdiff >>
rect -45 -215 225 -210
rect -45 -245 -30 -215
rect 210 -245 225 -215
rect -45 -250 225 -245
<< nsubdiff >>
rect -55 175 225 180
rect -55 145 -40 175
rect 210 145 225 175
rect -55 135 225 145
<< psubdiffcont >>
rect -30 -245 210 -215
<< nsubdiffcont >>
rect -40 145 210 175
<< poly >>
rect 0 80 15 95
rect 165 80 180 95
rect 0 -60 15 -15
rect -40 -65 15 -60
rect -40 -85 -30 -65
rect -10 -85 15 -65
rect -40 -90 15 -85
rect -115 -120 -100 -105
rect 0 -120 15 -90
rect 165 -35 180 -15
rect 165 -40 220 -35
rect 165 -60 190 -40
rect 210 -60 220 -40
rect 165 -65 220 -60
rect 165 -120 180 -65
rect 280 -120 295 -105
rect -115 -270 -100 -180
rect 0 -195 15 -180
rect 165 -195 180 -180
rect 280 -270 295 -180
rect -115 -285 295 -270
rect 50 -290 125 -285
rect 50 -315 60 -290
rect 115 -315 125 -290
rect 50 -320 125 -315
<< polycont >>
rect -30 -85 -10 -65
rect 190 -60 210 -40
rect 60 -315 115 -290
<< locali >>
rect -55 175 225 180
rect -55 145 -40 175
rect 210 145 225 175
rect -55 135 225 145
rect -30 75 -10 135
rect 190 75 215 135
rect -35 65 -5 75
rect -35 0 -30 65
rect -10 0 -5 65
rect -35 -10 -5 0
rect 20 65 50 75
rect 20 0 25 65
rect 45 0 50 65
rect 20 -40 50 0
rect 20 -60 25 -40
rect 45 -60 50 -40
rect -95 -65 0 -60
rect -95 -85 -30 -65
rect -10 -85 0 -65
rect -95 -90 0 -85
rect -250 -125 -120 -120
rect -250 -175 -240 -125
rect -215 -130 -120 -125
rect -215 -170 -145 -130
rect -125 -170 -120 -130
rect -215 -175 -120 -170
rect -250 -180 -120 -175
rect -95 -130 -65 -90
rect -95 -170 -90 -130
rect -70 -170 -65 -130
rect -95 -180 -65 -170
rect -35 -130 -5 -120
rect -35 -170 -30 -130
rect -10 -170 -5 -130
rect -35 -180 -5 -170
rect 20 -130 50 -60
rect 20 -170 25 -130
rect 45 -170 50 -130
rect 20 -180 50 -170
rect 130 65 160 75
rect 130 0 135 65
rect 155 0 160 65
rect 130 -90 160 0
rect 185 65 215 75
rect 185 0 190 65
rect 210 0 215 65
rect 185 -10 215 0
rect 180 -40 275 -35
rect 180 -60 190 -40
rect 210 -60 275 -40
rect 180 -65 275 -60
rect 130 -110 135 -90
rect 155 -110 160 -90
rect 130 -130 160 -110
rect 130 -170 135 -130
rect 155 -170 160 -130
rect 130 -180 160 -170
rect 185 -130 215 -120
rect 185 -170 190 -130
rect 210 -170 215 -130
rect 185 -180 215 -170
rect 245 -130 275 -65
rect 245 -170 250 -130
rect 270 -170 275 -130
rect 245 -180 275 -170
rect 300 -125 430 -120
rect 300 -130 395 -125
rect 300 -170 305 -130
rect 325 -170 395 -130
rect 300 -175 395 -170
rect 420 -175 430 -125
rect 300 -180 430 -175
rect -30 -210 -10 -180
rect 190 -210 210 -180
rect -45 -215 225 -210
rect -45 -245 -30 -215
rect 210 -245 225 -215
rect -45 -250 225 -245
rect 50 -290 125 -285
rect 50 -315 60 -290
rect 115 -315 125 -290
rect 50 -320 125 -315
<< viali >>
rect -40 145 210 175
rect 25 -60 45 -40
rect -240 -175 -215 -125
rect 135 -110 155 -90
rect 395 -175 420 -125
rect -30 -245 210 -215
<< metal1 >>
rect -55 175 225 180
rect -55 145 -40 175
rect 210 145 225 175
rect -55 135 225 145
rect -250 -125 -205 105
rect 20 -35 50 -30
rect 20 -40 210 -35
rect 20 -60 25 -40
rect 45 -60 210 -40
rect -40 -90 0 -60
rect 20 -65 210 -60
rect 20 -70 50 -65
rect 130 -90 160 -80
rect -40 -110 135 -90
rect 155 -110 160 -90
rect 130 -120 160 -110
rect -250 -175 -240 -125
rect -215 -175 -205 -125
rect -250 -250 -205 -175
rect 385 -125 430 105
rect 385 -175 395 -125
rect 420 -175 430 -125
rect -45 -215 225 -210
rect -45 -245 -30 -215
rect 210 -245 225 -215
rect -45 -250 225 -245
rect 385 -250 430 -175
rect 50 -340 125 -285
rect -175 -380 355 -340
<< via1 >>
rect -40 145 210 175
rect -30 -245 210 -215
<< metal2 >>
rect -180 175 375 180
rect -180 145 -40 175
rect 210 145 375 175
rect -180 135 375 145
rect -165 -215 345 -210
rect -165 -245 -30 -215
rect 210 -245 345 -215
rect -165 -250 345 -245
<< end >>
